library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ip is port
(
	pt	:	in std_logic_vector(1 TO 64);
	l0x	:	out std_logic_vector(1 TO 32);
	r0x	:	out std_logic_vector(1 TO 32)
);
end ip;

architecture behavior of ip is
begin
	l0x(1)<=pt(58);		l0x(2)<=pt(50);		l0x(3)<=pt(42);		l0x(4)<=pt(34);		l0x(5)<=pt(26);		l0x(6)<=pt(18);		l0x(7)<=pt(10);		l0x(8)<=pt(2);
	l0x(9)<=pt(60);		l0x(10)<=pt(52);	l0x(11)<=pt(44);	l0x(12)<=pt(36);	l0x(13)<=pt(28);	l0x(14)<=pt(20);	l0x(15)<=pt(12);	l0x(16)<=pt(4);
	l0x(17)<=pt(62);	l0x(18)<=pt(54);	l0x(19)<=pt(46);	l0x(20)<=pt(38);	l0x(21)<=pt(30);	l0x(22)<=pt(22);	l0x(23)<=pt(14);	l0x(24)<=pt(6);
	l0x(25)<=pt(64);	l0x(26)<=pt(56);	l0x(27)<=pt(48);	l0x(28)<=pt(40);	l0x(29)<=pt(32);	l0x(30)<=pt(24);	l0x(31)<=pt(16);	l0x(32)<=pt(8);

	r0x(1)<=pt(57);		r0x(2)<=pt(49);		r0x(3)<=pt(41);		r0x(4)<=pt(33);		r0x(5)<=pt(25);		r0x(6)<=pt(17);		r0x(7)<=pt(9);		r0x(8)<=pt(1);
	r0x(9)<=pt(59);		r0x(10)<=pt(51);	r0x(11)<=pt(43);	r0x(12)<=pt(35);	r0x(13)<=pt(27);	r0x(14)<=pt(19);	r0x(15)<=pt(11);	r0x(16)<=pt(3);
	r0x(17)<=pt(61);	r0x(18)<=pt(53);	r0x(19)<=pt(45);	r0x(20)<=pt(37);	r0x(21)<=pt(29);	r0x(22)<=pt(21);	r0x(23)<=pt(13);	r0x(24)<=pt(5);
	r0x(25)<=pt(63);	r0x(26)<=pt(55);	r0x(27)<=pt(47);	r0x(28)<=pt(39);	r0x(29)<=pt(31);	r0x(30)<=pt(23);	r0x(31)<=pt(15);	r0x(32)<=pt(7);
end behavior;
