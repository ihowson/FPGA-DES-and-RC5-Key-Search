library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fp is port
(      
	l,r	:	in	std_logic_vector(1 to 32);
	ct	:	out	std_logic_vector(1 to 64)
);
end fp;                                  

architecture behaviour of fp is
begin
	ct(1)<=r(8);	ct(2)<=l(8);	ct(3)<=r(16);	ct(4)<=l(16);	ct(5)<=r(24);	ct(6)<=l(24);	ct(7)<=r(32);	ct(8)<=l(32);
	ct(9)<=r(7);	ct(10)<=l(7);	ct(11)<=r(15);	ct(12)<=l(15);	ct(13)<=r(23);	ct(14)<=l(23);	ct(15)<=r(31);	ct(16)<=l(31);
	ct(17)<=r(6);	ct(18)<=l(6);	ct(19)<=r(14);	ct(20)<=l(14);	ct(21)<=r(22);	ct(22)<=l(22);	ct(23)<=r(30);	ct(24)<=l(30);
	ct(25)<=r(5);	ct(26)<=l(5);	ct(27)<=r(13);	ct(28)<=l(13);	ct(29)<=r(21);	ct(30)<=l(21);	ct(31)<=r(29);	ct(32)<=l(29);
	ct(33)<=r(4);	ct(34)<=l(4);	ct(35)<=r(12);	ct(36)<=l(12);	ct(37)<=r(20);	ct(38)<=l(20);	ct(39)<=r(28);	ct(40)<=l(28);
	ct(41)<=r(3);	ct(42)<=l(3);	ct(43)<=r(11);	ct(44)<=l(11);	ct(45)<=r(19);	ct(46)<=l(19);	ct(47)<=r(27);	ct(48)<=l(27);
	ct(49)<=r(2);	ct(50)<=l(2);	ct(51)<=r(10);	ct(52)<=l(10);	ct(53)<=r(18);	ct(54)<=l(18);	ct(55)<=r(26);	ct(56)<=l(26);
	ct(57)<=r(1);	ct(58)<=l(1);	ct(59)<=r(9);	ct(60)<=l(9);	ct(61)<=r(17);	ct(62)<=l(17);	ct(63)<=r(25);	ct(64)<=l(25);
end;
